library verilog;
use verilog.vl_types.all;
entity milestone1_tb is
end milestone1_tb;
